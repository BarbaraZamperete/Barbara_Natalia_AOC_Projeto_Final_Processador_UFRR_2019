LIBRARY ieee; 
USE ieee.std_logic_1164.all; 
USE ieee.numeric_std.all;  
USE ieee.std_logic_unsigned.all;

ENTITY ExtensorIS
	PORT(
		ENTRADA : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		ENTRADA2: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		SAIDA   : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		extend : IN STD_LOGIC
	);
	
END Extensor;

ARCHITECTURE BEHAVIOR OF Extensor  IS

BEGIN
 process(ENTRADA, ENTRADA2)
  begin
	if(extend = '1') then
			SAIDA <= ("00000") & ENTRADA;		
	end if;
	if(extend = '0') then
			SAIDA <= ("0000") & ENTRADA2;		
	end if;
 end process;
END BEHAVIOR;